`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/17/09 23:39:02
// Design Name: 
// Module Name: Shift
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`include "constant.v"

module Shift(
    input [16:0] state,
    input [5:0] r_dis4,
    input [5:0] r_dis3,
    input [5:0] r_dis2,
    input [5:0] r_dis1,
    input [5:0] dis_3,
    input [5:0] dis_2,
    input [5:0] dis_1,
    input clk,
    output reg [5:0] display0=`dis0,
    output reg [5:0] display1=`dis0,
    output reg [5:0] display2=`dis0,
    output reg [5:0] display3=`dis0,
    output reg [5:0] display4=`dis0,
    output reg [5:0] display5=`dis0,
    output reg [5:0] display6=`dis0,
    output reg [5:0] display7=`dis0
);
always@(posedge clk)begin
    case(state)
        `s1:begin
            display7<=`dis0;
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;
        end
        `s2:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;//0
        end
        `s3:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis1;//1
        end
        `s4:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis2;//2
        end
        `s5:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis3;//3
        end
        `s6:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis4;//4
        end
        `s7:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis5;//5
        end
        `s8:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis6;//6
        end
        `s9:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis7;//7
        end
        `s10:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis0;//0
        end
        `s11:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis1;//1
        end
        `s12:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis2;//2
        end
        `s13:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis3;//3
        end
        `s14:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis4;//4
        end
        `s15:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis5;//5
        end
        `s16:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis6;//6
        end
        `s17:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis13;//l
            display1<=`dis14;//o
            display0<=`dis7;//7
        end
        `s18:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis0;//0
        end
        `s19:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis1;//1
        end
        `s20:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis2;//2
        end
        `s21:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis3;//3
        end
        `s22:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis4;//4
        end
        `s23:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis5;//5
        end
        `s24:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis6;//6
        end
        `s25:begin
            display7<=`dis10;//F
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis15;//H
            display3<=`dis16;//i
            display2<=`dis17;//g
            display1<=`dis18;//h
            display0<=`dis7;//7
        end
        `s26:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;//0
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;
        end
        `s27:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;//0
        end
        `s28:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis1;//1
        end
        `s29:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis2;//2
        end
        `s30:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis3;//3
        end
        `s31:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis4;//4
        end
        `s32:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis5;//5
        end
        `s33:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis6;//6
        end
        `s34:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis1;//1
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis7;//7
        end
        `s35:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis2;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;//0
        end
        `s36:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis2;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis1;//1
        end
        `s37:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis2;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis2;//2
        end
        `s38:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis2;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis3;//3
        end
        `s39:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis2;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis4;//4
        end
        `s40:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis2;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis5;//5
        end
        `s41:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis2;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis6;//6
        end
        `s42:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;//2
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis7;//7
        end
        `s43:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;//0
        end
        `s44:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis1;//1
        end
        `s45:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis2;//2
        end
        `s46:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis3;//3
        end
        `s47:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis4;//4
        end
        `s48:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis5;//5
        end
        `s49:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis6;//6
        end
        `s50:begin
            display7<=`dis11;//A
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis3;//3
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis7;//7
        end
        `s51:begin//record
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=r_dis4;
            display3<=r_dis3;
            display2<=r_dis2;
            display1<=r_dis1;
            display0<=`dis0;//0
        end
        `s52:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis21;//c
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;//0
        end
        `s53:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis21;//c
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s54:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis21;//c
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s55:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis21;//c
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s56:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis21;//c
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s57:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis22;//d
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;//0
        end
        `s58:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis22;//d
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s59:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis22;//d
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s60:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis22;//d
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s61:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis22;//d
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s62:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis19;//E
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;//0
        end
        `s63:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis19;//E
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s64:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis19;//E
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s65:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis19;//E
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s66:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis19;//E
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s67:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis10;//F
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;//0
        end
        `s68:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis10;//F
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s69:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis10;//F
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s70:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis10;//F
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s71:begin
            display7<=`dis12;//S
            display6<=`dis0;
            display5<=`dis0;
            display4<=`dis10;//F
            display3<=dis_3;
            display2<=dis_2;
            display1<=dis_1;
            display0<=`dis0;
        end
        `s72:begin
            display7<=`dis20;//r
            display6<=`dis23;//e
            display5<=`dis21;//c
            display4<=`dis14;//o
            display3<=`dis20;//r
            display2<=`dis22;//d
            display1<=`dis0;
            display0<=`dis0;
        end
        `s73:begin
            display7<=`dis11;//A
            display6<=`dis22;//d
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;
        end
        `s74:begin
            display7<=`dis20;//r
            display6<=`dis22;//d
            display5<=`dis0;
            display4<=`dis0;
            display3<=`dis0;
            display2<=`dis0;
            display1<=`dis0;
            display0<=`dis0;
        end
    endcase
end
endmodule
