`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/12/22 22:20:20
// Design Name: 
// Module Name: pic
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`include "constant.v"
//This module is aim to generate the displayed image for VGA
module vga_pic(
input clk,
input rst_n,
input [2:0] mode,
input [2:0] select,//song select
input [9:0] pix_x,//x of the valid region
input [9:0] pix_y,//y of the valid region
output reg [11:0] pix_data//VGA display information
    );

reg [9:0] char_x;//Displays the legal area of the information
reg [9:0] char_y;
reg [9:0] char_a_x;
reg [9:0] char_a_y;

reg [255:0] char [63:0];//the area of the information for 4 characters
reg [511:0] cchar [63:0]; //the legal area of the information for 8 characters
reg [511:0] char_a[31:0];

always@(*) begin
if(((pix_x >= `aCHAR_B_H) && (pix_x < `aCHAR_B_H + `aCHAR_W)) && ((pix_y >= `aCHAR_B_V) && (pix_y < `aCHAR_B_V + `aCHAR_H))) begin
char_a_x = pix_x - `aCHAR_B_H;
char_a_y = pix_y - `aCHAR_B_V;
end else begin
char_a_x = 10'h3ff;
char_a_y = 10'h3ff;
end
end

always@ (*)  begin//Determines the display range of characters
case({mode, select})
`auto_s0, `auto_s1, `auto_s2: begin
if(((pix_x >= `cCHAR_B_H) && (pix_x < `cCHAR_B_H + `cCHAR_W)) && ((pix_y >= `cCHAR_B_V) && (pix_y < `cCHAR_B_V + `cCHAR_H))) begin
char_x = pix_x - `cCHAR_B_H;
char_y = pix_y - `cCHAR_B_V;
end else begin
char_x = 10'h3ff;
char_y = 10'h3ff;
end
end

default: begin
if(((pix_x >= `CHAR_B_H) && (pix_x < `CHAR_B_H + `CHAR_W)) && ((pix_y >= `CHAR_B_V) && (pix_y < `CHAR_B_V + `CHAR_H))) begin
char_x = pix_x - `CHAR_B_H;
char_y = pix_y - `CHAR_B_V;
end else begin
char_x = 10'h3ff;
char_y = 10'h3ff;
end
end

endcase
end

always@ (posedge clk)begin
char_a[0] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[1] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[2] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[3] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[4] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[5] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[6] <= 512'h000000000000000000000000000000000000000000000000000000000000000002000000000C0000000000000000000003006000000000000000000000060000;
char_a[7] <= 512'h0000000007C003C07FFC0000000000003000000000000000000000000000000006000000001800001FFFFF801FFFFF80020060000FFFFFC0000FFFE0000F0000;
char_a[8] <= 512'h0000000018300C30000C000000000000300000000000000000000000000000000600000000100000000600001000008006006000080000C07FCFFFE000198000;
char_a[9] <= 512'h00000000201818180018000000000000000000000000100000000000000000000600FFC03FFFFFE000060000100000800C3FFFC0080000C0060180000030C000;
char_a[10] <= 512'h00000000000830080010000000000000000000000000100000000000000000007FF880C0006000003FFFFFC010000080180060000FFFFFC00601800000E07000;
char_a[11] <= 512'h00C000000008200C0030000000000000000000000000100000000000000000007FF880C000C000002006004013FFFC8010C06000080000000601000001801800;
char_a[12] <= 512'h0FF81FC00008200C006033F833C007F0300007E007F0FF0000000000000000000C1080C00180000027E67E40100000802198618008FFFF800601000006000700;
char_a[13] <= 512'h1E183000001820040040340C3400180C300018180C0010000000000000000000081080C003FFFF0000060000100000807F18618008008000060300003FFFFDC0;
char_a[14] <= 512'h380020000010600400C038063800300630003008100010000000000000000000083080C007000300000600001000008002186180080080000603000060000040;
char_a[15] <= 512'h700020000060600400803002300020023000200C200010000000000000000000183080C00F00030007E67E0010FFF0800618618008FFFF800603FFC000000000;
char_a[16] <= 512'h7000300000C0600401803003300020023000200C200010000000000000000000182080C03B0003000000000010C030800C18618008C081800600008000000000;
char_a[17] <= 512'h70001C0003006004010030033000600330007FFC600010000000000000000000106080C063FFFF000FFFFF0010C030801818618008C081800600008000000000;
char_a[18] <= 512'h700003000C0020040300300330006003300060006000100000000000000000001C6080C0430003000806010010C03080309FFF80083FFE000600008007FFFE00;
char_a[19] <= 512'h700000C01800200C02003002300060033000600060001000000000000000000006C080C0030003000806010010C030803F806000080080000600008004000200;
char_a[20] <= 512'h7000004030003008060030023000200230002000200010000000000000000000038080C0030003000806010010C030800000600009FFFFC00600008004000200;
char_a[21] <= 512'h780000402000101804003806300030063000300030001000000000000000000001C080C003FFFF000FFFFF0010FFF080000060201900804007F0008004000200;
char_a[22] <= 512'h3C1800C06000183004003C0C3000180C30001808180018000000000000000000037080C003000300080601001000008000006020110084407F80008004000200;
char_a[23] <= 512'h1FF83F807FF807E00C0033F0300007F030000FF007F00F0000000000000000000E18FFC00300030008060100100000801FC06060313FFE406000018004000200;
char_a[24] <= 512'h03C0000000000000000030000000000030000000000000000000000000000000180880C003000300080601001000008070006060210000400000030007FFFE00;
char_a[25] <= 512'h0000000000000000000030000000000030000000000000000000000000000000700080C00300FE000FFFFF0010003F8000003FC0610009C00001FE0004000200;
char_a[26] <= 512'h00000000000000000000300000000000200000000000000000000000000000000000000003000000080001000000000000000000010006000000000004000200;
char_a[27] <= 512'h00000000000000000000300000000000600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[28] <= 512'h00000000000000000000300000000000C00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[29] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[30] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char_a[31] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end


always@ (posedge clk) begin
case(mode)
`mode_free ://free mode
begin
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h000000E000000000000000000000000000000000000000000000000000000000;
char[4] <= 256'h000000FC0000000000000000000000000008000003C000000000000000000000;
char[5] <= 256'h000000FE000000000000000000000000000F000003E00000000000F800000000;
char[6] <= 256'h000000FE000000000000001E00000000000F800003C00000000000781E000000;
char[7] <= 256'h000000FC000000000000001F800000000007003C03C00000000000780FC00000;
char[8] <= 256'h000000F8000000000000000F800000000007001E038000000000003807E00000;
char[9] <= 256'h000001F0000000000000000F800000000007000E038400000000003803E00000;
char[10] <= 256'h000001E0000000000000000F800000000007000E03FF00000000003800E00000;
char[11] <= 256'h000001E0000000000000000F800000000007000E3FFE00000000001800600000;
char[12] <= 256'h000003C00000000000000007000000000007000FFF8000000000001800000000;
char[13] <= 256'h00000380000000000000000700000000000703FFC60000000000001C00000000;
char[14] <= 256'h000007807E0000000000000700000000000301F7040000000000001C00000000;
char[15] <= 256'h0000070FFF800000000000070000000000030003040000000000001C00000000;
char[16] <= 256'h0001FFFFFFC00000000000070000000000032003080000000000000C78000000;
char[17] <= 256'h0003FFFC1FE0000000000007000000000003F801006000000000000FFC000000;
char[18] <= 256'h0001FC001FF0000000000007001F0000001FF00007F000000000003FF8000000;
char[19] <= 256'h0001F0000FE000000000000707FFC00000FFC003FCFC0000000001FFC0000000;
char[20] <= 256'h0001F0000FE0000000040007FFFFE0000FFF007E007C000000001FFE00000000;
char[21] <= 256'h0001F0000FC00000000780FFF807F0000FCF0070007800000003FFE700000000;
char[22] <= 256'h0001F0000FC000000007FFFF0003F000000F0030007000000003FC0700000000;
char[23] <= 256'h0000F0000FC000000003F0070003E000000F0039F8F000000000000300000000;
char[24] <= 256'h0000F0000FC000000003C0070003E000001F003FF0E000000000000380000000;
char[25] <= 256'h0000F01F07C000000003C0070003C000001FC01800E000000000000380000000;
char[26] <= 256'h0000F3FF87C000000003C0070003C000003BF01801C000000000000180000000;
char[27] <= 256'h0000FFFF87C000000001C0070003C000003B78180FC0000000000001C0000000;
char[28] <= 256'h0000FFFC07C000000001C0070003C0000077381BFF800000000001C1C0000000;
char[29] <= 256'h0000FE0007C000000001C0070003C0000077180FC100000000000FF0E0000000;
char[30] <= 256'h0000F00007C000000001C0071E03C00000E70008E00000000000FFE0E0000000;
char[31] <= 256'h0000F00007C000000001C007FF03800000C7000070000000000FFF0060000000;
char[32] <= 256'h0000F00007C000000001C7FFFF03800001C70000601F80000007FC0070000000;
char[33] <= 256'h0000F03F07C000000001C7FFF0078000038700006FFFC00000001E0078000000;
char[34] <= 256'h0000FFFF87C000000001C3E7000780000307000FFFFFE00000001E0038000000;
char[35] <= 256'h0000FFFF87C000000000E0070007800006071FFFE000000000000E001C000000;
char[36] <= 256'h0001FFFE07C000000000E007000780000C070FF8E000000000000C001C000000;
char[37] <= 256'h0001F00007C000000000E0070007800018070100F000000000000C060E000000;
char[38] <= 256'h0001F00007C000000000E0070007800010070001D800000000000CFC0F000000;
char[39] <= 256'h0001F00007C000000000E0070007800020070001CC00000000000FF007000000;
char[40] <= 256'h0001F00007C000000000E00700070000000700018E00000000003F8007801000;
char[41] <= 256'h0001F00007C000000000E0070007000000070003870000000001FC0003C01000;
char[42] <= 256'h0001F01FCFC000000000E0073F8F0000000E000703800000000FF00001E01000;
char[43] <= 256'h0001FFFFFFC000000000607FFFCF0000000E000E03E0000001FF800000F01000;
char[44] <= 256'h0001FFFFFFC0000000006FFFFFFF0000000E001E01F0000001FE000000F83000;
char[45] <= 256'h0001FC007FC0000000007FE0007F0000000E003800FC000000F80000007E3000;
char[46] <= 256'h0001E0003FC0000000006000003E0000000E00F0007F000000000000003F7000;
char[47] <= 256'h0000E0003F80000000006000003E0000000603C0003FC00000000000001FF000;
char[48] <= 256'h0000E0001F80000000002000003E000000060C00001FF00000000000000FF000;
char[49] <= 256'h000000001F80000000000000001C000000000000000FF000000000000003F800;
char[50] <= 256'h000000000F00000000000000001C00000000000000000000000000000001F800;
char[51] <= 256'h000000000F000000000000000018000000000000000000000000000000007800;
char[52] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end
`mode_auto ://auto
begin
    if(select == `sel_s1)begin
cchar[0] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[1] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[2] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[3] <= 512'h000000E00000000000000000000000000000000000000000000001E0000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[4] <= 512'h000000FC0000000000000000000000000000000700000000000000F0000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[5] <= 512'h000000FE00000000000000000000000000000003C0000000000000F0000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[6] <= 512'h000000FE00000000000000000080000000000003E0000000000000E00000000000000000000000000000008000000000000000000F000000000000000F000000;
cchar[7] <= 512'h000000FC000000000000000000F0000000000001F0000000000000E0000000000000000000000000000000F00000000000000001FFC0000000000001FFC00000;
cchar[8] <= 512'h000000F8000000000000000000F80000003C0000F0000000000000E1F800000000000000000000000000007C000000000000007FE7F000000000007FE7F00000;
cchar[9] <= 512'h000001F0000000000000000000F80000001F000060000000000001FFFC00000000000000000000000000003E000000000001FFF003F800000001FFF003F80000;
cchar[10] <= 512'h000001E0000000000000000000F00000001F80002018000000003FFFF000000000000000000000000000003E000000000001FC0003F800000001FC0003F80000;
cchar[11] <= 512'h000001E0000000000000000000F00000000F800001FE000000003FF80000000000000000000000000000003C000000000000F00003E000000000F00003E00000;
cchar[12] <= 512'h000003C0000000000000000000F00000000780001FFF8000000001C00000000000000000000000000000003C000000000000780103E000000000780103E00000;
cchar[13] <= 512'h00000380000000000000000000F0000000038C01FF1FC000000001C00000000000000000000000000000003C000000000000781FC3C000000000781FC3C00000;
cchar[14] <= 512'h000007807E0000000000000000E0000000000C7FE01FC000000001C00000000000000000000000000000003C00000000000039FF87800000000039FF87800000;
cchar[15] <= 512'h0000070FFF800000000000FC00E0000000001FF8001E00000000018FF000000000000000000000000000001C0000000000003FF80780000000003FF807800000;
cchar[16] <= 512'h0001FFFFFFC0000000003FFE00E0000000001C0000180000000003FFF000000000000000000000000000001C0000000000001C000700000000001C0007000000;
cchar[17] <= 512'h0003FFFC1FE000000001FFE000E0000000003C00002000000000FFFE0000000000000000000000000000001C0000000000001C000F00000000001C000F000000;
cchar[18] <= 512'h0001FC001FF0000000007C0000E0E000000038003C00000000007F000000000000000000000000000000001C0000000000000C000E00000000000C000E000000;
cchar[19] <= 512'h0001F0000FE000000000000001E3F80000007801FC000000000003000000000000000000000000000000001C0000000000000C03FE00000000000C03FE000000;
cchar[20] <= 512'h0001F0000FE000000000000001FFFC000300701FF0000000000007001C00000000000000000000000000001C0000000000000EFFFC00000000000EFFFC000000;
cchar[21] <= 512'h0001F0000FC00000000000001FF87E0007E0703FC000000000000707FF00000000000000000000000000001C00000000000007F808000000000007F808000000;
cchar[22] <= 512'h0001F0000FC00000000000007FC07C0003F0200700000000000007FFFF00000000000000000000000000001C0180000000000638000000000000063800000000;
cchar[23] <= 512'h0000F0000FC000000000000639C03C0001F000038180000000007FFF0000000000000000000000000004001C01F000000000001E000000000000001E00000000;
cchar[24] <= 512'h0000F0000FC000000000007F83C0380000F000038FE00000003FFF8600000000000E0000000000000004001C00F800000000001E000000000000001E00000000;
cchar[25] <= 512'h0000F01F07C0000000000FFF0380380000200003FFF80000001FEC0300000000001F800000000000000C001C007E00000000C01E000000000000C01E00000000;
cchar[26] <= 512'h0000F3FF87C000000003FFC00380780000001C3FC1F8000000001C0180000000003F800000000000000C001C003E00000000F01C000000000000F01C00000000;
cchar[27] <= 512'h0000FFFF87C0000001FFF0000380780000000FFB80F0000000001C00C0000000003FC00000000000001C001C003F00000000F81C000000000000F81C00000000;
cchar[28] <= 512'h0000FFFC07C0000000FF1C000780700000000E0380F000000000380070000000003FC00000000000001C001C001F80000001F01C7F8000000001F01C7F800000;
cchar[29] <= 512'h0000FE0007C0000000001C00070070000001070381E000000000380038000000003F800000000000003C001C000F80000001E01FFF8000000001E01FFF800000;
cchar[30] <= 512'h0000F00007C0000000003C000700700000020703F9E00000000070061E000000001F800000000000003C001C000FC0000003C3FFFC0000000003C3FFFC000000;
cchar[31] <= 512'h0000F00007C00000000038000F0070000002031FF1C000000000E03F1F000000000E000000000000007C001C0007C0000007FFFF000000000007FFFF00000000;
cchar[32] <= 512'h0000F00007C00000000030600E0070000006033F81C000000001E7FE0F800000000000000000000000F8001C0003C000000F3F9C00000000000F3F9C00000000;
cchar[33] <= 512'h0000F03F07C00000000070700E007000000C030381C000000003CFF007E00000000000000000000000F8001C00038000001E001C00000000001E001C00000000;
cchar[34] <= 512'h0000FFFF87C00000000060381E00F000000C030303800000000381C003F80000000000000000000001F0001C000180000038001C000000000038001C00000000;
cchar[35] <= 512'h0000FFFF87C000000000C07C1C00E0000018030303800000000F01C001FF0000000000000000000001F0001C000000000070001C000000000070001C00000000;
cchar[36] <= 512'h0001FFFE07C000000000C3DE1C00E00000380183FF000000001E01C1E0FFE000000000000000000000E0001C000000000080001C7C0000000080001C7C000000;
cchar[37] <= 512'h0001F00007C000000001DF0E3800E000003801FFFF000000003801FFF87FF800000000000000000000C0001C000000000000001FFF0000000000001FFF000000;
cchar[38] <= 512'h0001F00007C000000003FC0E3800E000007001F00200000000701FFFF800000000000000000000000000001C00000000000003FFFF000000000003FFFF000000;
cchar[39] <= 512'h0001F00007C00000000FF0067001E00000F000800000000001C3FFF80000000000000000000000000000001C0000000000003FFF0000000000003FFF00000000;
cchar[40] <= 512'h0001F00007C00000000FC0007001C00001E000400000000007007B800000000000000000000000000000003C0000000000000F9C0000000000000F9C00000000;
cchar[41] <= 512'h0001F00007C00000000F0000E001C00003E00070100000000000038000000000001F0000000000000000003C000000000000001C000000000000001C00000000;
cchar[42] <= 512'h0001F01FCFC0000000060001E003C00003E000F80E0000000000038000000000003F80000000000000001C3C000000000000001C000000000000001C00000000;
cchar[43] <= 512'h0001FFFFFFC0000000000001C003C00001E000F8078000000000070600000000003FC00000000000000007FC000000000000001C000000000000001C00000000;
cchar[44] <= 512'h0001FFFFFFC00000000000038107800001C001F003E000000000070380000000003FC00000000000000003FC000000000000001C001F80000000001C001F8000;
cchar[45] <= 512'h0001FC007FC000000000000701EF800000C003C001F0000000000E01E0000000003FC00000000000000001F8000000000000001C7FFFE0000000001C7FFFE000;
cchar[46] <= 512'h0001E0003FC000000000000E00FF00000040078000F8000000001C01F8000000003F800000000000000001F800000000000001FFFFFFF000000001FFFFFFF000;
cchar[47] <= 512'h0000E0003F8000000000001C007F000000000E00007C000000007800FC000000001F000000000000000000F000000000000FFFFFFFFFF800000FFFFFFFFFF800;
cchar[48] <= 512'h0000E0001F80000000000038007E000000001C00007C00000001F0007C000000000000000000000000000070000000000FFFFFE0000000000FFFFFE000000000;
cchar[49] <= 512'h000000001F80000000000070003C000000003000003C0000000780003E0000000000000000000000000000200000000007FFE0000000000007FFE00000000000;
cchar[50] <= 512'h000000000F000000000000C0003800000000C00000180000000000003E0000000000000000000000000000000000000001E000000000000001E0000000000000;
cchar[51] <= 512'h000000000F00000000000100001000000000000000000000000000001E0000000000000000000000000000000000000000000000000000000000000000000000;
cchar[52] <= 512'h000000000000000000000000000000000000000000000000000000000C0000000000000000000000000000000000000000000000000000000000000000000000;
cchar[53] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[54] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[55] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[56] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[57] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[58] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[59] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[60] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[61] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[62] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[63] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end else if(select == `sel_s2)begin
cchar[0] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[1] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[2] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[3] <= 512'h000000E00000000000000000000000000000000000000000000001E0000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[4] <= 512'h000000FC0000000000000000000000000000000700000000000000F0000000000000000000000000000000018000000000000000000000000000000000000000;
cchar[5] <= 512'h000000FE00000000000000000000000000000003C0000000000000F000000000000000000000000000000001E000000000000000700000000000000000000000;
cchar[6] <= 512'h000000FE00000000000000000080000000000003E0000000000000E000000000000000000000000000000001F0000000000000007C0000000000000000000000;
cchar[7] <= 512'h000000FC000000000000000000F0000000000001F0000000000000E000000000000000000000000000000001F000000000000000FE0000000000000000000000;
cchar[8] <= 512'h000000F8000000000000000000F80000003C0000F0000000000000E1F8000000000000000000000000000001E000000000000003FF0000000000000000030000;
cchar[9] <= 512'h000001F0000000000000000000F80000001F000060000000000001FFFC000000000000000000000000000001E00000000000000FFF00000000000000007FE000;
cchar[10] <= 512'h000001E0000000000000000000F00000001F80002018000000003FFFF0000000000000000000000000000001C00000000000007F80000000000000001FFFE000;
cchar[11] <= 512'h000001E0000000000000000000F00000000F800001FE000000003FF800000000000000000000000000000003C0000000000183F8000000000018001FFFFC0000;
cchar[12] <= 512'h000003C0000000000000000000F00000000780001FFF8000000001C000000000000000000000000000000003800000000000FF8000000000001E000FF8000000;
cchar[13] <= 512'h00000380000000000000000000F0000000038C01FF1FC000000001C000000000000000000000000000000003800000000000F80000000000001F0E001C000000;
cchar[14] <= 512'h000007807E0000000000000000E0000000000C7FE01FC000000001C000000000000000000000000000000007000000000000E00000000000001E0F803C000000;
cchar[15] <= 512'h0000070FFF800000000000FC00E0000000001FF8001E00000000018FF0000000000000000000000000000007000000000000E07000000000001E07C038000000;
cchar[16] <= 512'h0001FFFFFFC0000000003FFE00E0000000001C0000180000000003FFF000000000000000000000000000780F00C000000000E03E00000000001C03E030000000;
cchar[17] <= 512'h0003FFFC1FE000000001FFE000E0000000003C00002000000000FFFE0000000000000000000000000003FC0E03F000000000E03F00000000003C01E060700000;
cchar[18] <= 512'h0001FC001FF0000000007C0000E0E000000038003C00000000007F0000000000000000000000000003FFFC0E1FFC00000000E01E00000000003800E047FC0000;
cchar[19] <= 512'h0001F0000FE000000000000001E3F80000007801FC0000000000030000000000000000000000000007FC7C1DFFFE00000000E01E000000000038006FFFBF0000;
cchar[20] <= 512'h0001F0000FE000000000000001FFFC000300701FF0000000000007001C000000000000000000000001C0781FE0FC00000000C01C000000000070000FC00F0000;
cchar[21] <= 512'h0001F0000FC00000000000001FF87E0007E0703FC000000000000707FF00000000000000000000000000703800F000000000C01C000000000071C006000F0000;
cchar[22] <= 512'h0001F0000FC00000000000007FC07C0003F0200700000000000007FFFF00000000000000000000000000707001C000000001C01C07F0000000E1E006000E0000;
cchar[23] <= 512'h0000F0000FC000000000000639C03C0001F000038180000000007FFF00000000000000000000000000007060018000000001C01FFFF8000000C1F0060C0E0000;
cchar[24] <= 512'h0000F0000FC000000000007F83C0380000F000038FE00000003FFF8600000000000E0000000000000000E0C4010000000003C0FFFFF0000001C1E0060F0E0000;
cchar[25] <= 512'h0000F01F07C0000000000FFF0380380000200003FFF80000001FEC0300000000001F80000000000000C0E087000000000007FFFFC00000000381C0060F0E0000;
cchar[26] <= 512'h0000F3FF87C000000003FFC00380780000001C3FC1F8000000001C0180000000003F8000000000000070E007C00000000007FFDC00000000030180060E0E0000;
cchar[27] <= 512'h0000FFFF87C0000001FFF0000380780000000FFB80F0000000001C00C0000000003FC000000000000038E007800000000007F01C00000000060380060E0E0000;
cchar[28] <= 512'h0000FFFC07C0000000FF1C000780700000000E0380F000000000380070000000003FC00000000000001DC007800000000007001C000000000C0300060E0E0000;
cchar[29] <= 512'h0000FE0007C0000000001C00070070000001070381E000000000380038000000003F800000000000000FC007800000000000001C00000000100700060E0E0000;
cchar[30] <= 512'h0000F00007C0000000003C000700700000020703F9E00000000070061E000000001F800000000000000FC007800000000000001C00000000000618060E0E0000;
cchar[31] <= 512'h0000F00007C00000000038000F0070000002031FF1C000000000E03F1F000000000E00000000000000078007800000000000001C00000000000E1E060E0E0000;
cchar[32] <= 512'h0000F00007C00000000030600E0070000006033F81C000000001E7FE0F80000000000000000000000003C007800000000000001C00000000000C0F0E0E0E0000;
cchar[33] <= 512'h0000F03F07C00000000070700E007000000C030381C000000003CFF007E0000000000000000000000007E007C00000000000001C00000000001C0F8E0E0E0000;
cchar[34] <= 512'h0000FFFF87C00000000060381E00F000000C030303800000000381C003F8000000000000000000000007F007C00000000001801C1E0000000018078E0E0E0000;
cchar[35] <= 512'h0000FFFF87C000000000C07C1C00E0000018030303800000000F01C001FF00000000000000000000000EF807600000000003801C0FC00000003FFFCE1C0E0000;
cchar[36] <= 512'h0001FFFE07C000000000C3DE1C00E00000380183FF000000001E01C1E0FFE0000000000000000000001E780E700000000003801C07F00000007FE3CC1C0E0000;
cchar[37] <= 512'h0001F00007C000000001DF0E3800E000003801FFFF000000003801FFF87FF8000000000000000000001C7C0E300000000007801C03F8000001FF01841C0E0000;
cchar[38] <= 512'h0001F00007C000000003FC0E3800E000007001F00200000000701FFFF8000000000000000000000000383C0C38000000000F801C01FC000001FC00001C0E0000;
cchar[39] <= 512'h0001F00007C00000000FF0067001E00000F000800000000001C3FFF800000000000000000000000000781C1C1C000000000F001C00FE000001F0000039840000;
cchar[40] <= 512'h0001F00007C00000000FC0007001C00001E000400000000007007B8000000000000000000000000000701C1C0E000000001F001C007E000000C0000078E00000;
cchar[41] <= 512'h0001F00007C00000000F0000E001C00003E00070100000000000038000000000001F00000000000000E008380F000000003E001C003F00000000000070780000;
cchar[42] <= 512'h0001F01FCFC0000000060001E003C00003E000F80E0000000000038000000000003F80000000000001C0007007800000003E001C001F000000000000F07C0000;
cchar[43] <= 512'h0001FFFFFFC0000000000001C003C00001E000F8078000000000070600000000003FC000000000000380007007C00000003C001C000F000000000001E03E0000;
cchar[44] <= 512'h0001FFFFFFC00000000000038107800001C001F003E000000000070380000000003FC00000000000060000E003F000000038001C0007000000000003C01F0000;
cchar[45] <= 512'h0001FC007FC000000000000701EF800000C003C001F0000000000E01E0000000003FC000000000000C0001C003F800000000073C0000000000000007800F0000;
cchar[46] <= 512'h0001E0003FC000000000000E00FF00000040078000F8000000001C01F8000000003F8000000000000000070001FE0000000003FC000000000000000E000F0000;
cchar[47] <= 512'h0000E0003F8000000000001C007F000000000E00007C000000007800FC000000001F00000000000000000E0001FFC000000001FC000000000000003800070000;
cchar[48] <= 512'h0000E0001F80000000000038007E000000001C00007C00000001F0007C00000000000000000000000000300000FFF000000000FC00000000000000E000030000;
cchar[49] <= 512'h000000001F80000000000070003C000000003000003C0000000780003E000000000000000000000000000000001F800000000078000000000000000000010000;
cchar[50] <= 512'h000000000F000000000000C0003800000000C00000180000000000003E0000000000000000000000000000000000000000000078000000000000000000000000;
cchar[51] <= 512'h000000000F00000000000100001000000000000000000000000000001E0000000000000000000000000000000000000000000030000000000000000000000000;
cchar[52] <= 512'h000000000000000000000000000000000000000000000000000000000C0000000000000000000000000000000000000000000000000000000000000000000000;
cchar[53] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[54] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[55] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[56] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[57] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[58] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[59] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[60] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[61] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[62] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[63] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end else if(select == `sel_s3)begin
cchar[0] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[1] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[2] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[3] <= 512'h000000E00000000000000000000000000000000000000000000001E0000000000000000000000000000000F00000000000000000000000000000003000000000;
cchar[4] <= 512'h000000FC0000000000000000000000000000000700000000000000F0000000000000000000000000000000F80000000000000000000000000000003C00000000;
cchar[5] <= 512'h000000FE00000000000000000000000000000003C0000000000000F00000000000000000000000000000007C0000000000000000000000000000003E00000000;
cchar[6] <= 512'h000000FE00000000000000000080000000000003E0000000000000E00000000000000000000000000000003C000000000000C0000C0000000000001F00000000;
cchar[7] <= 512'h000000FC000000000000000000F0000000000001F0000000000000E00000000000000000000000000000001C000000000000F0000F8000000000000F00000000;
cchar[8] <= 512'h000000F8000000000000000000F80000003C0000F0000000000000E1F800000000000000000000000000000003F000000000F8001FC000000000000600000000;
cchar[9] <= 512'h000001F0000000000000000000F80000001F000060000000000001FFFC000000000000000000000000000003FFF800000000F8001FC00000000000000FC00000;
cchar[10] <= 512'h000001E0000000000000000000F00000001F80002018000000003FFFF00000000000000000000000000001FFFFFC00000000F0003F00000000000001FFC00000;
cchar[11] <= 512'h000001E0000000000000000000F00000000F800001FE000000003FF8000000000000000000000000007FFFFFC00000000001E0007C0000000000001FFF800000;
cchar[12] <= 512'h000003C0000000000000000000F00000000780001FFF8000000001C0000000000000000000000000003FFF00000000000001E001F0000000000003FFF8000000;
cchar[13] <= 512'h00000380000000000000000000F0000000038C01FF1FC000000001C0000000000000000000000000001F0000000000000001C003C000000000007FFE60000000;
cchar[14] <= 512'h000007807E0000000000000000E0000000000C7FE01FC000000001C000000000000000000000000000000000000000000003C007C000000000003FC078000000;
cchar[15] <= 512'h0000070FFF800000000000FC00E0000000001FF8001E00000000018FF0000000000000000000000000000003E00000000003801DE00000000000000078000000;
cchar[16] <= 512'h0001FFFFFFC0000000003FFE00E0000000001C0000180000000003FFF000000000000000000000000000007FF0000000000781F0E00000000000000078000000;
cchar[17] <= 512'h0003FFFC1FE000000001FFE000E0000000003C00002000000000FFFE00000000000000000000000000007FF9F0000000000700E0E000000000000E0070000000;
cchar[18] <= 512'h0001FC001FF0000000007C0000E0E000000038003C00000000007F0000000000000000000000000000003C01F0000000000F00E0E000000000000700E0000000;
cchar[19] <= 512'h0001F0000FE000000000000001E3F80000007801FC0000000000030000000000000000000000000000003C01E0000000000E00E07000000000000780C0000000;
cchar[20] <= 512'h0001F0000FE000000000000001FFFC000300701FF0000000000007001C000000000000000000000000001C01C0000000001E00E0701C000000000380C0000000;
cchar[21] <= 512'h0001F0000FC00000000000001FF87E0007E0703FC000000000000707FF000000000000000000000000001C0180000000001C0060707E00000000038180000000;
cchar[22] <= 512'h0001F0000FC00000000000007FC07C0003F0200700000000000007FFFF000000000000000000000000000C1FC0000000003E006071FC00000000018183FFE000;
cchar[23] <= 512'h0000F0000FC000000000000639C03C0001F000038180000000007FFF00000000000000000000000000000FFF80000000003F00603FF0000000000007FFFFF800;
cchar[24] <= 512'h0000F0000FC000000000007F83C0380000F000038FE00000003FFF8600000000000E00000000000000000F8000000000007300603FC00000000003FFFFFFF800;
cchar[25] <= 512'h0000F01F07C0000000000FFF0380380000200003FFF80000001FEC0300000000001F800000000000000004000060000000E38060FE0000000003FFFC00000000;
cchar[26] <= 512'h0000F3FF87C000000003FFC00380780000001C3FC1F8000000001C0180000000003F8000000000000000000003F8000000E38067F800000007FFFC0000000000;
cchar[27] <= 512'h0000FFFF87C0000001FFF0000380780000000FFB80F0000000001C00C0000000003FC0000000000000000003FFFE000001C380679C00000007FF800000000000;
cchar[28] <= 512'h0000FFFC07C0000000FF1C000780700000000E0380F000000000380070000000003FC00000000000008007FFFFFF0000038380601C00000003F0000000000000;
cchar[29] <= 512'h0000FE0007C0000000001C00070070000001070381E000000000380038000000003F80000000000000FFFFE0003F0000070380600E0000000000000078000000;
cchar[30] <= 512'h0000F00007C0000000003C000700700000020703F9E00000000070061E000000001F80000000000000FFE000001F00000C0380E00E00000000000003FE000000;
cchar[31] <= 512'h0000F00007C00000000038000F0070000002031FF1C000000000E03F1F000000000E00000000000000700000001E0000080380E00F000000000000FFFF000000;
cchar[32] <= 512'h0000F00007C00000000030600E0070000006033F81C000000001E7FE0F800000000000000000000000700003001E0000000300E00700000000003FF01F800000;
cchar[33] <= 512'h0000F03F07C00000000070700E007000000C030381C000000003CFF007E0000000000000000000000070003FC01C0000000300E04780000000001C001F000000;
cchar[34] <= 512'h0000FFFF87C00000000060381E00F000000C030303800000000381C003F8000000000000000000000070FFFFE01C0000000300E08380000000001C000F000000;
cchar[35] <= 512'h0000FFFF87C000000000C07C1C00E0000018030303800000000F01C001FF0000000000000000000000707E03E01C0000000300E303C0000000001C000E000000;
cchar[36] <= 512'h0001FFFE07C000000000C3DE1C00E00000380183FF000000001E01C1E0FFE000000000000000000000707803C01C0000000300E701C0000000001C000E000000;
cchar[37] <= 512'h0001F00007C000000001DF0E3800E000003801FFFF000000003801FFF87FF800000000000000000000703803801C0000000300EE01E0100000001C070E000000;
cchar[38] <= 512'h0001F00007C000000003FC0E3800E000007001F00200000000701FFFF8000000000000000000000000703803001C0000000700FC00F0100000001DFF8E000000;
cchar[39] <= 512'h0001F00007C00000000FF0067001E00000F000800000000001C3FFF800000000000000000000000000703803001C0000000701F80070100000001FFE0E000000;
cchar[40] <= 512'h0001F00007C00000000FC0007001C00001E000400000000007007B80000000000000000000000000007019FF801C0000000703F1F078100000001C000E000000;
cchar[41] <= 512'h0001F00007C00000000F0000E001C00003E00070100000000000038000000000001F00000000000000701FFF001C0000000703E0FC3C100000001C000E000000;
cchar[42] <= 512'h0001F01FCFC0000000060001E003C00003E000F80E0000000000038000000000003F80000000000000701800001C0000000703C07C1E300000001C000E000000;
cchar[43] <= 512'h0001FFFFFFC0000000000001C003C00001E000F8078000000000070600000000003FC0000000000000700800001C0000000F03C03C0FB00000001C000E000000;
cchar[44] <= 512'h0001FFFFFFC00000000000038107800001C001F003E000000000070380000000003FC0000000000000700000003C0000000F01801C07F00000001C001E000000;
cchar[45] <= 512'h0001FC007FC000000000000701EF800000C003C001F0000000000E01E0000000003FC0000000000000700000003C0000000F00000007F00000001C3FDE000000;
cchar[46] <= 512'h0001E0003FC000000000000E00FF00000040078000F8000000001C01F8000000003F80000000000000700000387C0000000F00000003F80000001FFFFE000000;
cchar[47] <= 512'h0000E0003F8000000000001C007F000000000E00007C000000007800FC000000001F000000000000007000000FFC0000000E00000001F80000001F003E000000;
cchar[48] <= 512'h0000E0001F80000000000038007E000000001C00007C00000001F0007C00000000000000000000000020000007F80000000600000000780000000C003E000000;
cchar[49] <= 512'h000000001F80000000000070003C000000003000003C0000000780003E00000000000000000000000020000003F80000000600000000380000000C001C000000;
cchar[50] <= 512'h000000000F000000000000C0003800000000C00000180000000000003E00000000000000000000000000000001F000000000000000000000000000001C000000;
cchar[51] <= 512'h000000000F00000000000100001000000000000000000000000000001E00000000000000000000000000000001E0000000000000000000000000000008000000;
cchar[52] <= 512'h000000000000000000000000000000000000000000000000000000000C00000000000000000000000000000000C0000000000000000000000000000000000000;
cchar[53] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[54] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[55] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[56] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[57] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[58] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[59] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[60] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[61] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[62] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
cchar[63] <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end else begin//direct display �Զ�����
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h000000E00000000000000000000000000000000000000000000001E000000000;
char[4] <= 256'h000000FC0000000000000000000000000000000700000000000000F000000000;
char[5] <= 256'h000000FE00000000000000000000000000000003C0000000000000F000000000;
char[6] <= 256'h000000FE00000000000000000080000000000003E0000000000000E000000000;
char[7] <= 256'h000000FC000000000000000000F0000000000001F0000000000000E000000000;
char[8] <= 256'h000000F8000000000000000000F80000003C0000F0000000000000E1F8000000;
char[9] <= 256'h000001F0000000000000000000F80000001F000060000000000001FFFC000000;
char[10] <= 256'h000001E0000000000000000000F00000001F80002018000000003FFFF0000000;
char[11] <= 256'h000001E0000000000000000000F00000000F800001FE000000003FF800000000;
char[12] <= 256'h000003C0000000000000000000F00000000780001FFF8000000001C000000000;
char[13] <= 256'h00000380000000000000000000F0000000038C01FF1FC000000001C000000000;
char[14] <= 256'h000007807E0000000000000000E0000000000C7FE01FC000000001C000000000;
char[15] <= 256'h0000070FFF800000000000FC00E0000000001FF8001E00000000018FF0000000;
char[16] <= 256'h0001FFFFFFC0000000003FFE00E0000000001C0000180000000003FFF0000000;
char[17] <= 256'h0003FFFC1FE000000001FFE000E0000000003C00002000000000FFFE00000000;
char[18] <= 256'h0001FC001FF0000000007C0000E0E000000038003C00000000007F0000000000;
char[19] <= 256'h0001F0000FE000000000000001E3F80000007801FC0000000000030000000000;
char[20] <= 256'h0001F0000FE000000000000001FFFC000300701FF0000000000007001C000000;
char[21] <= 256'h0001F0000FC00000000000001FF87E0007E0703FC000000000000707FF000000;
char[22] <= 256'h0001F0000FC00000000000007FC07C0003F0200700000000000007FFFF000000;
char[23] <= 256'h0000F0000FC000000000000639C03C0001F000038180000000007FFF00000000;
char[24] <= 256'h0000F0000FC000000000007F83C0380000F000038FE00000003FFF8600000000;
char[25] <= 256'h0000F01F07C0000000000FFF0380380000200003FFF80000001FEC0300000000;
char[26] <= 256'h0000F3FF87C000000003FFC00380780000001C3FC1F8000000001C0180000000;
char[27] <= 256'h0000FFFF87C0000001FFF0000380780000000FFB80F0000000001C00C0000000;
char[28] <= 256'h0000FFFC07C0000000FF1C000780700000000E0380F000000000380070000000;
char[29] <= 256'h0000FE0007C0000000001C00070070000001070381E000000000380038000000;
char[30] <= 256'h0000F00007C0000000003C000700700000020703F9E00000000070061E000000;
char[31] <= 256'h0000F00007C00000000038000F0070000002031FF1C000000000E03F1F000000;
char[32] <= 256'h0000F00007C00000000030600E0070000006033F81C000000001E7FE0F800000;
char[33] <= 256'h0000F03F07C00000000070700E007000000C030381C000000003CFF007E00000;
char[34] <= 256'h0000FFFF87C00000000060381E00F000000C030303800000000381C003F80000;
char[35] <= 256'h0000FFFF87C000000000C07C1C00E0000018030303800000000F01C001FF0000;
char[36] <= 256'h0001FFFE07C000000000C3DE1C00E00000380183FF000000001E01C1E0FFE000;
char[37] <= 256'h0001F00007C000000001DF0E3800E000003801FFFF000000003801FFF87FF800;
char[38] <= 256'h0001F00007C000000003FC0E3800E000007001F00200000000701FFFF8000000;
char[39] <= 256'h0001F00007C00000000FF0067001E00000F000800000000001C3FFF800000000;
char[40] <= 256'h0001F00007C00000000FC0007001C00001E000400000000007007B8000000000;
char[41] <= 256'h0001F00007C00000000F0000E001C00003E00070100000000000038000000000;
char[42] <= 256'h0001F01FCFC0000000060001E003C00003E000F80E0000000000038000000000;
char[43] <= 256'h0001FFFFFFC0000000000001C003C00001E000F8078000000000070600000000;
char[44] <= 256'h0001FFFFFFC00000000000038107800001C001F003E000000000070380000000;
char[45] <= 256'h0001FC007FC000000000000701EF800000C003C001F0000000000E01E0000000;
char[46] <= 256'h0001E0003FC000000000000E00FF00000040078000F8000000001C01F8000000;
char[47] <= 256'h0000E0003F8000000000001C007F000000000E00007C000000007800FC000000;
char[48] <= 256'h0000E0001F80000000000038007E000000001C00007C00000001F0007C000000;
char[49] <= 256'h000000001F80000000000070003C000000003000003C0000000780003E000000;
char[50] <= 256'h000000000F000000000000C0003800000000C00000180000000000003E000000;
char[51] <= 256'h000000000F00000000000100001000000000000000000000000000001E000000;
char[52] <= 256'h000000000000000000000000000000000000000000000000000000000C000000;
char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end
end
`mode_study://study 
begin
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h000000001E000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h000000001F800000000000000000000000000000000000000000000000000000;
char[4] <= 256'h000000001FC0000000000000000000000008000003C000000000000000000000;
char[5] <= 256'h000000E01FC000000000000000000000000F000003E00000000000F800000000;
char[6] <= 256'h0001C0F81F8000000000000000000000000F800003C00000000000781E000000;
char[7] <= 256'h0001F07C1F00000000000000000000000007003C03C00000000000780FC00000;
char[8] <= 256'h0000F87C3E00000000000000000000000007001E038000000000003807E00000;
char[9] <= 256'h0000FC7E3E0000000000000000E000000007000E038400000000003803E00000;
char[10] <= 256'h0000FC3E3C0000000000000007F800000007000E03FF00000000003800E00000;
char[11] <= 256'h00007C3C7800000000000000FFFE00000007000E3FFE00000000001800600000;
char[12] <= 256'h00003C1C78000000000001FFFFFF00000007000FFF8000000000001800000000;
char[13] <= 256'h00003C00F000000000003FFF003F0000000703FFC60000000000001C00000000;
char[14] <= 256'h00001800E0FF000000001FC0003E0000000301F7040000000000001C00000000;
char[15] <= 256'h00000001FFFF800000000000001E000000030003040000000000001C00000000;
char[16] <= 256'h0030003FFFFFC00000000000001E000000032003080000000000000C78000000;
char[17] <= 256'h00783FFFF01FE00000000000001C00000003F801006000000000000FFC000000;
char[18] <= 256'h007FFFF0001FF00000000000001C0000001FF00007F000000000003FF8000000;
char[19] <= 256'h007FF800003FF00000000000001C000000FFC003FCFC0000000001FFC0000000;
char[20] <= 256'h00F80000003F800000000200001C00000FFF007E007C000000001FFE00000000;
char[21] <= 256'h00F80007007C0000000003C0001C00000FCF0070007800000003FFE700000000;
char[22] <= 256'h01F0007FC0700000000003F0001C0000000F0030007000000003FC0700000000;
char[23] <= 256'h01F03FFFE0E00000000001F8001C0000000F0039F8F000000000000300000000;
char[24] <= 256'h03F1FFE7F0000000000000F8001C0000001F003FF0E000000000000380000000;
char[25] <= 256'h03E0FF07F000000000000078001C0000001FC01800E000000000000380000000;
char[26] <= 256'h03E0700FC000000000000038001C0000003BF01801C000000000000180000000;
char[27] <= 256'h01C0000F0000000000000018001C0000003B78180FC0000000000001C0000000;
char[28] <= 256'h0000001E0000000000000000001C00000077381BFF800000000001C1C0000000;
char[29] <= 256'h000000F80000000000000000181C00000077180FC100000000000FF0E0000000;
char[30] <= 256'h0000007801F8000000000000601C000000E70008E00000000000FFE0E0000000;
char[31] <= 256'h0000007FFFFF000000000001C01C000000C7000070000000000FFF0060000000;
char[32] <= 256'h0000007FFFFF000000000007801C000001C70000601F80000007FC0070000000;
char[33] <= 256'h00007FFFFFFF80000000001E003C0000038700006FFFC00000001E0078000000;
char[34] <= 256'h03FFFFFE000300000000007C003C00000307000FFFFFE00000001E0038000000;
char[35] <= 256'h07FFFF1E00000000000001F8003C000006071FFFE000000000000E001C000000;
char[36] <= 256'h03FFC01F00000000000007E0003C00000C070FF8E000000000000C001C000000;
char[37] <= 256'h00F0001F0000000000001FC0003C000018070100F000000000000C060E000000;
char[38] <= 256'h0000001F000000000003FF000038000010070001D800000000000CFC0F000000;
char[39] <= 256'h0000001F000000000003FE000038000020070001CC00000000000FF007000000;
char[40] <= 256'h0000001F000000000001FC0000780000000700018E00000000003F8007801000;
char[41] <= 256'h0000001F000000000000F8000078000000070003870000000001FC0003C01000;
char[42] <= 256'h0000001F000000000000700000780000000E000703800000000FF00001E01000;
char[43] <= 256'h0000001F000000000000000000F80000000E000E03E0000001FF800000F01000;
char[44] <= 256'h0000001F000000000000000180F00000000E001E01F0000001FE000000F83000;
char[45] <= 256'h0000001F00000000000000007FF00000000E003800FC000000F80000007E3000;
char[46] <= 256'h0000003F00000000000000003FF00000000E00F0007F000000000000003F7000;
char[47] <= 256'h00001F7E00000000000000001FE00000000603C0003FC00000000000001FF000;
char[48] <= 256'h00000FFE00000000000000000FC0000000060C00001FF00000000000000FF000;
char[49] <= 256'h000007FE00000000000000000FC0000000000000000FF000000000000003F800;
char[50] <= 256'h000003FC0000000000000000078000000000000000000000000000000001F800;
char[51] <= 256'h000001F800000000000000000600000000000000000000000000000000007800;
char[52] <= 256'h000000F000000000000000000000000000000000000000000000000000000000;
char[53] <= 256'h000000E000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end
`mode_record: begin
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h0000000000000000000000000000000000000000000000000000003000000000;
char[4] <= 256'h0000000000000000000000000000000000000000000000000000003C00000000;
char[5] <= 256'h0000000000000000000000000000000000000000000000000000003E00000000;
char[6] <= 256'h0000000000000000000100001000000000000000FC0000000000001F00000000;
char[7] <= 256'h00000000000000000001C0001C0000000000000FFE0000000000000F00000000;
char[8] <= 256'h0000000003C000000001F0001E000000000003FFFF0000000000000600000000;
char[9] <= 256'h00000000FFE000000000F0001F0000000003FFF03F000000000000000FC00000;
char[10] <= 256'h0000003FFFF000000000F0001E0000000000FC003E00000000000001FFC00000;
char[11] <= 256'h00007FFFFF8000000000E0001E000000000000003C0000000000001FFF800000;
char[12] <= 256'h0007FFFFC00000000000E0003C000000000000003C000000000003FFF8000000;
char[13] <= 256'h0001FF81E00000000000E0003800000000000007B800000000007FFE60000000;
char[14] <= 256'h00001E00F00000000000E00038000000000001FFF800000000003FC078000000;
char[15] <= 256'h00000E00F00000000000C0007000000000001FFF700000000000000078000000;
char[16] <= 256'h00000F00F00000000000C0007000000000000780700000000000000078000000;
char[17] <= 256'h00000F00F00000000001C00060000000000000006000000000000E0070000000;
char[18] <= 256'h00000F00E00000000001C000E0700000000000006078000000000700E0000000;
char[19] <= 256'h00000E00E00000000001C000C07C0000000000007FFE000000000780C0000000;
char[20] <= 256'h00000E00E000000000018601C03F00000000001FFFFE000000000380C0000000;
char[21] <= 256'h00000E00E007C00000018381801F800000003FFFFE0600000000038180000000;
char[22] <= 256'h00000E00EFFFF000000183C3000FC00000FFFFF0000000000000018183FFE000;
char[23] <= 256'h00000E0FFFFFF00000018387003FC00000FFF8700000000000000007FFFFF800;
char[24] <= 256'h0000FFFFFFFC000000038F8F1FFFE000003E007802000000000003FFFFFFF800;
char[25] <= 256'h0FFFFFFF600000000003FF1FFF81E00000000038038000000003FFFC00000000;
char[26] <= 256'h07FFFE0060000000003FC71FF80040000000003803C0000007FFFC0000000000;
char[27] <= 256'h03F80E00600000001FFF071F800000000000003803E0000007FF800000000000;
char[28] <= 256'h00000E00600000001FF3060C000000000000003807C0000003F0000000000000;
char[29] <= 256'h00000C00600000000F870E00000000000003F03E0E0000000000000078000000;
char[30] <= 256'h00000C007000000000070E00000000000001F0371C00000000000003FE000000;
char[31] <= 256'h00001C007000000000060E00000000000000F033B0000000000000FFFF000000;
char[32] <= 256'h00001C007000000000060C000000000000007039C000000000003FF01F800000;
char[33] <= 256'h00001C007000000000071C00007E000000000038E000000000001C001F000000;
char[34] <= 256'h000018007000000000039C0007FF8000000000387000000000001C000F000000;
char[35] <= 256'h00003800700000000001F80FFFFFC000000000383800000000001C000E000000;
char[36] <= 256'h00003800700000000000F80FE00F8000000002383E00000000001C000E000000;
char[37] <= 256'h000070007000000000007007000F0000000004381F00000000001C070E000000;
char[38] <= 256'h000070007000000000007807000F0000000018380F80000000001DFF8E000000;
char[39] <= 256'h0000E000700000000000FC07000E00000000703807E0000000001FFE0E000000;
char[40] <= 256'h0000C000700000000001DE07001E00000000E03803F8000000001C000E000000;
char[41] <= 256'h0001C0007000000000038F03001C00000003C03801FF000000001C000E000000;
char[42] <= 256'h000380007000000000070F03001C0000003F803800FFE00000001C000E000000;
char[43] <= 256'h0007000060000000001E0703007C0000007F0038007FF80000001C000E000000;
char[44] <= 256'h000600006000000000380303BFFE0000003F00380008000000001C001E000000;
char[45] <= 256'h000C00006000000000700201FFE00000000E00380000000000001C3FDE000000;
char[46] <= 256'h00100000600000000180000180000000000007780000000000001FFFFE000000;
char[47] <= 256'h00000000600000000000000100000000000003F80000000000001F003E000000;
char[48] <= 256'h00000000600000000000000000000000000001F80000000000000C003E000000;
char[49] <= 256'h00000000600000000000000000000000000001F00000000000000C001C000000;
char[50] <= 256'h00000000600000000000000000000000000000F000000000000000001C000000;
char[51] <= 256'h0000000020000000000000000000000000000060000000000000000008000000;
char[52] <= 256'h0000000000000000000000000000000000000040000000000000000000000000;
char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end
`mode_read: begin
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h0000000000000000000000000000000000000000000000000000003000000000;
char[4] <= 256'h0000000000000000000000001C00000000000000000000000000003C00000000;
char[5] <= 256'h0006000000000000000000001F00000000000000000000000000003E00000000;
char[6] <= 256'h000380000E000000000000001F00000000000000FC0000000000001F00000000;
char[7] <= 256'h0003C0001F0000000000F0001F0000000000000FFE0000000000000F00000000;
char[8] <= 256'h0003C0003F80000000007C001E000000000003FFFF0000000000000600000000;
char[9] <= 256'h0003C0007C00000000003E001E0000000003FFF03F000000000000000FC00000;
char[10] <= 256'h00038000E0E0000000003F003C0000000000FC003E00000000000001FFC00000;
char[11] <= 256'h00018003C0F8000000001F003C000000000000003C0000000000001FFF800000;
char[12] <= 256'h0001800CE0F0000000000F0038000000000000003C000000000003FFF8000000;
char[13] <= 256'h0001804071C00000000000003800000000000007B800000000007FFE60000000;
char[14] <= 256'h00018070718000000000000070000000000001FFF800000000003FC078000000;
char[15] <= 256'h0001807062000000000000007000000000001FFF700000000000000078000000;
char[16] <= 256'h000180386000000000000000E000000000000780700000000000000078000000;
char[17] <= 256'h000180186070000000000000E0020000000000006000000000000E0070000000;
char[18] <= 256'h0001F00067FC0000000003F0C01F8000000000006078000000000700E0000000;
char[19] <= 256'h0001F8007FFC000000003FE1C0FF8000000000007FFE000000000780C0000000;
char[20] <= 256'h000FF00FFF0000000007FE018FFE00000000001FFFFE000000000380C0000000;
char[21] <= 256'h007F83FFF000000001FFE003FFF0000000003FFFFE0600000000038180000000;
char[22] <= 256'h03FF81F9FC0000001FFF00037F00000000FFFFF0000000000000018183FFE000;
char[23] <= 256'h01E18003EE00000007E1C0070300000000FFF8700000000000000007FFFFF800;
char[24] <= 256'h00018007678000000301E00E03C00000003E007802000000000003FFFFFFF800;
char[25] <= 256'h0001900761C000000001E00C03C0000000000038038000000003FFFC00000000;
char[26] <= 256'h0001E00E60F000000001C010038000000000003803C0000007FFFC0000000000;
char[27] <= 256'h0001C01C607C00000001C000038000000000003803E0000007FF800000000000;
char[28] <= 256'h00038038603F00000003FF00038000000000003807C0000003F0000000000000;
char[29] <= 256'h00078070E01FE00000039F8C070000000003F03E0E0000000000000078000000;
char[30] <= 256'h001D80E0E00FFC00000787C6070000000001F0371C00000000000003FE000000;
char[31] <= 256'h003981C06007F000000707C3070000000000F033B0000000000000FFFF000000;
char[32] <= 256'h00F1830060F00000000E07818600000000007039C000000000003FF01F800000;
char[33] <= 256'h01E186001FFC0000000E0781CE00000000000038E000000000001C001F000000;
char[34] <= 256'h07818007F83E0000001C0700EE000000000000387000000000001C000F000000;
char[35] <= 256'h3F0183FE603C0000001C07007C000000000000383800000000001C000E000000;
char[36] <= 256'h3E0181C0603C0000003807007C000000000002383E00000000001C000E000000;
char[37] <= 256'h1C0181C060380000007007003C000000000004381F00000000001C070E000000;
char[38] <= 256'h000180E07E38000000600E007C000000000018380F80000000001DFF8E000000;
char[39] <= 256'h000180E3FE38000000C00E00FE0000000000703807E0000000001FFE0E000000;
char[40] <= 256'h000380E7E038000001800E01EF0000000000E03803F8000000001C000E000000;
char[41] <= 256'h000380E06038000003001C03C78000000003C03801FF000000001C000E000000;
char[42] <= 256'h000380606038000006083C0783C00000003F803800FFE00000001C000E000000;
char[43] <= 256'h00638060607800000C06781E01F00000007F0038007FF80000001C000E000000;
char[44] <= 256'h003F80606F7000001003F8F801F80000003F00380008000000001C001E000000;
char[45] <= 256'h001F8067FFF000000003F00000FE0000000E00380000000000001C3FDE000000;
char[46] <= 256'h000F007F80F000000001F000007FC000000007780000000000001FFFFE000000;
char[47] <= 256'h00070030007000000001E000003FF800000003F80000000000001F003E000000;
char[48] <= 256'h00060020006000000000C000001FFC00000001F80000000000000C003E000000;
char[49] <= 256'h00020000006000000000000000000000000001F00000000000000C001C000000;
char[50] <= 256'h00000000000000000000000000000000000000F000000000000000001C000000;
char[51] <= 256'h0000000000000000000000000000000000000060000000000000000008000000;
char[52] <= 256'h0000000000000000000000000000000000000040000000000000000000000000;
char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end
`mode_adjust:begin
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h0000000000000000000040000000000000000000000000000000000000000000;
char[4] <= 256'h0000000000000000000078003000000000000000000000000000000000000000;
char[5] <= 256'h0007000000000000000038003C00000000038000000000000000000000000000;
char[6] <= 256'h001FE000003F8000000038003E0000000003E00180000000000200003C000000;
char[7] <= 256'h001FF00007FFC000000038003C0000000001E001E0000000000380001E000000;
char[8] <= 256'h000FF9E7FFFFE000000038003C0000000001E000F80000000003C0001E000000;
char[9] <= 256'h0003F9FFFF0FF00000003800380000000001C000F80000000003C0001E000000;
char[10] <= 256'h0001F8FF3E07F00000003FE0700000000001C0007C000000000780000E000000;
char[11] <= 256'h000020F83F07E0000003FF80700C00000001C0003C000000000700000E000000;
char[12] <= 256'h000000F83E07E000000FF800607E00000001C0001C000000000700000E000000;
char[13] <= 256'h000000783E07C00000003000E1FC00000001C00008000000000600000E7C0000;
char[14] <= 256'h000000783E07C00000003000DFF000000001C00000100000000E00000FFE0000;
char[15] <= 256'h000000783FE7C000000033F9FF0000000001C000007C0000000E1C00FFBE0000;
char[16] <= 256'h0000007BFFF7C00000007FF9838000000001C04007FF0000000CFE03FE3C0000;
char[17] <= 256'h0000007BFFE7C000007FF0F3038000000001DC603F1F8000001FFC000E1CE000;
char[18] <= 256'h00078078FE07C000003030E3038000000001FE63F01F0000001F80700E3FF000;
char[19] <= 256'h001FE0783E07C000003830E5870000000003F8FF003C0000003801F80EFFE000;
char[20] <= 256'h007FE0783E07C000001830E8C7000000001FC0E000300000003007F81FF80000;
char[21] <= 256'h1FFFE0783FFFC00000183FE06E00000001FFC1E00040000000700037FE380000;
char[22] <= 256'h1FFFC07FFFFFC000001FF8003E00000001F9C1C0C000000000600073EE380000;
char[23] <= 256'h0F87C07FFFFFC000001870001E0000000001C1C0F000000000C0F0600E300000;
char[24] <= 256'h000780FBF007C0000008F8001E0000000001C980F000000001C3F0600FF80000;
char[25] <= 256'h000780F80007C0000000FF803F8000000001D180F0000000019FE0603FF00000;
char[26] <= 256'h000780F80007C0000001F7C073C000000001E000E0000000031F00C3FE000000;
char[27] <= 256'h000F80F007E7C0000003B1C0E1F000000001E000C1000000070700C1CE000000;
char[28] <= 256'h000F80F7FFFFC000000730E380FE00000001C000C38FF000060701C00E700000;
char[29] <= 256'h000F00FFFFFFC000000C700E007FE0000003C001CFFFF8000C0701800FF80000;
char[30] <= 256'h000F00F7E1FFC00000387000003FF000000FC003FFFFF8001807FB81FFF00000;
char[31] <= 256'h000F00F7C1F7C00000707001F80F0000001FC3FFE3800000100FF3F3FE000000;
char[32] <= 256'h000F01F3C1E7C00000E0203FF8000000003DFFFB03800000207FC3F80E000000;
char[33] <= 256'h000F0DE3C1E7C00003800FFF800000000079DE030700000003FF00380E3C0000;
char[34] <= 256'h000F3DE3C1C7C00004001FF80000000001F1C0070700000000E600300FFE0000;
char[35] <= 256'h000FF9E3FFE7C0000000003C0000000003E1C0060F000000000600307FF80000;
char[36] <= 256'h001FF3E1FFE7C0000000003C000000000FC1C00F0E00000000060037FC000000;
char[37] <= 256'h001FE3C1FE07C00000000038000000003F81C007DE00000000060071CC000000;
char[38] <= 256'h001FC3C1C007C00000004038180000001F01C001FC00000000060F600C000000;
char[39] <= 256'h003F83C08007C00000007039FC0000000601C0003E000000000603E00C000000;
char[40] <= 256'h003F87800007C0000000783FE00000000001C0007FC00000000610E00C000000;
char[41] <= 256'h003F07800007C00000007838000000000001C000F7E00000000660F80C000000;
char[42] <= 256'h003E0F000007C00000003038000000000021C001E3F800000007C1DE0C000000;
char[43] <= 256'h003C0F0003EFC0000000303800000000001FC003C0FC0000000F818F84000000;
char[44] <= 256'h001C1E0003FFC0000000303800000000001FC007007E0000000F8383F8000000;
char[45] <= 256'h00001C0000FFC0000000303800000000000F801E003E0000001F0700FE000000;
char[46] <= 256'h00003800007FC00000003038FFF8000000078078001F0000001E0C007FC00000;
char[47] <= 256'h00007800003FC000000031FFFFFE0000000781E0000F0000001C18001FFFF000;
char[48] <= 256'h00007000001F80000007FFFFE0FE000000030700000200000000000007FFF800;
char[49] <= 256'h00000000000F000001FFFE000000000000030000000000000000000001FFC000;
char[50] <= 256'h00000000000E000000FE000000000000000000000000000000000000007E0000;
char[51] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[52] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end
default:begin
end
endcase
end

always@ (posedge clk, negedge rst_n) begin//Stored characters with data transmitted to the display
if(!rst_n)
pix_data <= `BLACK;
else begin
case({mode, select})
`auto_s1,`auto_s2,`auto_s0: begin//While playing three songs
if(((pix_x >= `cCHAR_B_H - 1) && (pix_x < `cCHAR_B_H + `cCHAR_W - 1)) 
                                 && ((pix_y >= `cCHAR_B_V) && (pix_y < `cCHAR_B_V + `cCHAR_H)) 
                                 && (cchar[char_y][511-char_x] == 1'b1))//Need to reverse
pix_data <= `WHITE;
else if(((pix_x >= `aCHAR_B_H - 1) && (pix_x < `aCHAR_B_H + `aCHAR_W - 1)) 
                                 && ((pix_y >= `aCHAR_B_V) && (pix_y < `aCHAR_B_V + `aCHAR_H)) 
                                 && (char_a[char_a_y][511-char_a_x] == 1'b1))//Need to reverse)
pix_data <= `BULE;
else
pix_data <= `BLACK;
end

default: begin
if(((pix_x >= `CHAR_B_H - 1) && (pix_x < `CHAR_B_H + `CHAR_W - 1)) 
                                 && ((pix_y >= `CHAR_B_V) && (pix_y < `CHAR_B_V + `CHAR_H)) 
                                 && (char[char_y][255-char_x] == 1'b1))//Need to reverse
pix_data <= `WHITE;
else if(((pix_x >= `aCHAR_B_H - 1) && (pix_x < `aCHAR_B_H + `aCHAR_W - 1)) 
                                 && ((pix_y >= `aCHAR_B_V) && (pix_y < `aCHAR_B_V + `aCHAR_H)) 
                                 && (char_a[char_a_y][511-char_a_x] == 1'b1))//Need to reverse)
pix_data <= `BULE;
else
pix_data <= `BLACK;
end
endcase
end
end
endmodule
